class cfg;
    // Integer fields with default values
    int latency = 1;
    int amount = 100;

endclass
