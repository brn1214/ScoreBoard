// TODO: create transaction class

    // class transaction;
    // ..
    // enclass

// Class must containt single-bit bit fields:
// signal_in and signal_out
class transaction;
    // Single-bit fields
    bit X1;
    bit X2;
	bit X3;
	bit Y1;



endclass
