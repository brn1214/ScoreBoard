// TODO: create interface

    // interface inv_if(input logic clk);
    // ..
    // endinterface

// Interface must contain single-bit logic fields:
// signal_in and signal_out

interface inv_if(input logic clk);
    // Single-bit logic fields
    logic X1;
    logic X2;	  
	logic X3;  
	logic Y1;
																   
endinterface
